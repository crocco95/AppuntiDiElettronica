-- libraries
library IEEE;
use IEE.std_logic_1164.all;

-- entity
entity esercizio_2 is
	port(
		X1, X0: in std_logic;
		CLK, RST: in std_logic;
		Q1, Q0: out std_logic
	);
end esercizio_2;

-- architecture
architecture esercizio_2_architecture of esercizio_2 is

end esercizio_2_architecture